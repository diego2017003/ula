LIBRARY ieee;
use ieee.std_logic_1164.all;
ENTITY MULTIPLEXADOR1BIT IS 
	PORT(
		Em1,Em2,Em3,Em4,Em5,Em6:IN STD_LOGIC;
		S0,S1,S2,S3:IN STD_LOGIC;
		Saida:OUT STD_LOGIC);
END MULTIPLEXADOR1BIT;
ARCHITECTURE mux1BIT OF MULTIPLEXADOR1BIT IS
SIGNAL i1,i2,i3,i4,i5,i6:STD_LOGIC;
BEGIN
i1<=(Em1)AND(NOT(s3))AND(NOT(s2))AND(NOT(s1))AND(NOT(s0));	
i2<=(Em2)AND(NOT(s3))AND(NOT(s2))AND(NOT(s1))AND((s0));
i3<=(Em3)AND(NOT(s3))AND(NOT(s2))AND((s1))AND(NOT(s0));
i4<=(Em4)AND(NOT(s3))AND(NOT(s2))AND((s1))AND((s0));
i5<=(Em5)AND(NOT(s3))AND((s2))AND(NOT(s1))AND(NOT(s0));
i6<=(Em6)AND(NOT(s3))AND((s2))AND(NOT(s1))AND((s0));
Saida<=(i1)OR(i2)OR(i3)OR(i4)OR(i5)OR(i6);
END mux1BIT;