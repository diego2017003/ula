LIBRARY ieee;
use ieee.std_logic_1164.all;
ENTITY SUBTRACAOC2 IS 
	PORT(
		SE1,SE2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		SUBOut:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		SignOut:OUT STD_LOGIC);
END SUBTRACAOC2;
ARCHITECTURE subtraic2 OF SUBTRACAOC2 IS
COMPONENT SOMA8BITS
	PORT(Carryin:IN BIT;
		X1,X2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		Sout:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	Carryout:OUT STD_LOGIC);
END COMPONENT;
COMPONENT INVERSOR
	PORT(
		E:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		nE:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;
SIGNAL INV:STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	INVERTEE2:INVERSOR PORT MAP(E=>SE2,nE=>INV);
	subtracao:SOMA8BITS PORT MAP(Carryin=>'1',X1=>SE1,X2=>INV,Sout=>SUBOut,Carryout=>SignOut);
END subtraic2;