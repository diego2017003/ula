LIBRARY ieee;
use ieee.std_logic_1164.all;
ENTITY COMPARADOR8BITS IS 
	PORT(
		SE81,SE82:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		SE8q,SM8t,SL8t:OUT STD_LOGIC);
END COMPARADOR8BITS;
ARCHITECTURE compara8BITs OF COMPARADOR8BITS IS
COMPONENT COMPARADOR1BIT 
PORT(
		SE1,SE2,SoEq,SoMt,SoLt:IN STD_LOGIC;
		SEq,SMt,SLt:OUT STD_LOGIC);
END COMPONENT;
SIGNAL S1:STD_LOGIC_VECTOR(23 DOWNTO 0);
BEGIN
	C:COMPARADOR1BIT PORT MAP(SE1=>SE81(7),SE2=>SE82(7),SoEq=>'1',SoMt=>'0',SoLt=>'0',SEq=>S1(0),SMt=>S1(1),SLt=>S1(2));
	C2:COMPARADOR1BIT PORT MAP(SE1=>SE81(6),SE2=>SE82(6),SoEq=>S1(0),SoMt=>S1(1),SoLt=>S1(2),SEq=>S1(3),SMt=>S1(4),SLt=>S1(5));
	C3:COMPARADOR1BIT PORT MAP(SE1=>SE81(5),SE2=>SE82(5),SoEq=>S1(3),SoMt=>S1(4),SoLt=>S1(5),SEq=>S1(6),SMt=>S1(7),SLt=>S1(8));
	C4:COMPARADOR1BIT PORT MAP(SE1=>SE81(4),SE2=>SE82(4),SoEq=>S1(6),SoMt=>S1(7),SoLt=>S1(8),SEq=>S1(9),SMt=>S1(10),SLt=>S1(11));
	C5:COMPARADOR1BIT PORT MAP(SE1=>SE81(3),SE2=>SE82(3),SoEq=>S1(9),SoMt=>S1(10),SoLt=>S1(11),SEq=>S1(12),SMt=>S1(13),SLt=>S1(14));
	C6:COMPARADOR1BIT PORT MAP(SE1=>SE81(2),SE2=>SE82(2),SoEq=>S1(12),SoMt=>S1(13),SoLt=>S1(14),SEq=>S1(15),SMt=>S1(16),SLt=>S1(17));
	C7:COMPARADOR1BIT PORT MAP(SE1=>SE81(1),SE2=>SE82(1),SoEq=>S1(15),SoMt=>S1(16),SoLt=>S1(17),SEq=>S1(18),SMt=>S1(19),SLt=>S1(20));
	C8:COMPARADOR1BIT PORT MAP(SE1=>SE81(0),SE2=>SE82(0),SoEq=>S1(18),SoMt=>S1(19),SoLt=>S1(20),SEq=>S1(21),SMt=>S1(22),SLt=>S1(23));

	SE8q<=S1(21);
	SM8t<=S1(22);
	SL8t<=S1(23);
END compara8BITs;